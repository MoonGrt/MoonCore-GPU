`timescale 1ns / 1ps

module Drv_MIPI (
    input wire clk,  // ʱ��
    input wire rstn  // ��λ���͵�ƽ��Ч

);



endmodule
